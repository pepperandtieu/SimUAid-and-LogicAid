�d d        d    ��  Cor3�   �����   v���                       ��  Cinput�   �����   ����0 0 A�   ����        ��   �����   ����1 1 Q2'�   ����        ��   }����   }���0 0 Q3�   ����         ��  Coutput�   �����   ����1 1                  ��  Cnand2  ����W  p���                       �  ����  ����1 1 S1'�   ����        �  }���  }���1 1                   �W  ����G  ����0 0 Q1W  ����        	��   �����   ����                       ��   �����   ����0 0 A�   ����        ��   �����   ����0 0 Q1�   ����         ��   �����   ����1 1                  ��  Cor2�   �����   s���                       ��   �����   ����0 0 B�   ����        ��   �����   ����0 0 Q2�   ����         ��   �����   ����0 0 R3'�   ����        	�  ����X  ����                       �  ����  ����1 1                  �  ����  ����1 1                   �W  ����I  ����0 0 Q3W  ����        ��  Cnand3  ����X  s���                       �  ����  ����0 0                  �  ����  ����0 0                  �  y���  y���1 1 R  ����         �W  ����I  ����1 1 Q3'W  ����        �  D���W  "���                       �  >���  >���0 0                  �  3���  3���1 1 Q3'�   <���        �  (���  (���1 1 R  ,���         �W  3���G  3���1 1 Q1'W  B���        	��  ����!  u���                       ��  �����  ����0 0 B�  ����        ��  �����  ����1 1 Q3'�  ����         �   ����  ����1 1 S2'!  ����        	�N  �����  p���                       �N  ����]  ����1 1                  �N  }���]  }���1 1                   ��  �����  ����0 0 Q2�  ����        	�N  �����  ����                       �N  ����]  ����1 1                  �N  ����]  ����1 1                   ��  �����  ����0 0 Z�  ����        	��  ����   q���                       ��  �����  ����0 0 A�  ����        ��  ����  ���1 1 Q2'�  ����         �   ����  ����1 1                  �N  E����  #���                       �N  ?���]  ?���0 0                  �N  4���]  4���1 1                  �N  )���]  )���1 1 RB  1���         ��  4����  4���1 1 Q2'�  3���        ��  ����   ����                       ��  �����  ����0 0 A�  ����        ��  �����  ����1 1 Q1'�  ����        ��  �����  ����1 1 Q3'�  ����         �   ����  ����1 1                  ��  F���  #���                       ��  9����  9���0 0 A�  D���        ��  /����  /���1 1 Q3'�  6���         �  4���  4���1 1 R2'  C���        ��  Cinput_signal   o���Q   ^���                         �Q   f���E   f���0 0                   ��  Csignal    0 G�   1 G�   0 G�   1 G�   0 G�#   1 G�-   0 ��  Cswitch   ����O   ����O   ����i   ���� R     �   ����.   ����1 Z                  �   ����.   ����0 Z                   �O   ����A   ����1 1 RO   ����        D�   ���S   ����                         �S   ���E   ���0 0                   G�    0 G�
   1 G�2   0 ��  Cprobe�  �����  �����  �����  ����  Z     ��  �����  ����0 0 Z�  ����          Y�n  �����  ����f  �����  ����  Q1     �x  ����x  ����0 0 Q1f  ����          Y��  �����  �����  �����  ����  Q2     ��  �����  ����0 0 Q2�  ����          Y�p  	����  ����l  ����  ���  Q3     �z  ����z  ����0 0 Q3l  ���          Y�W   ����k   f���d   ����}   ����  A     ��  Cpina   f���a   t���0 0 Ad   ����          Y�Z   #���n   ���g   5����   #���  B     c�d   ���d   ���0 0 Bg   5���           ��  Cnet1  ��  Csegment�   ����  ����i��   �����   ����i�  ����  ����    g�0 	 i��  T����  ����i�W  ����W  ����i�x  ����W  ����i��   T����  T���i�  >���  >���i��   >���  >���i��   T����   >���i��  ����x  ����i�x  ����x  ���� " ]    g�0  i��   ����  ����i��   �����   ����i�  ����  ����    g�1  i��   �����   ����i�  ����  ����i�v  �����   ����i�W  ����W  ����i�v  ����W  ����i�v  ����v  ����i�  �����   ����  # ( > B    g�0  i�  �����   ����i��   �����   ����i�  ����  ����i��  �����   ����i�W  ����W  ����i�W  ����W  ����i��  �����  ����i�z  ����W  ����i��  ����z  ����i�z  ����z  ����i�z  ����z  ����i�z  ����z  ����  a    g�1  i�   ����N  ����i�   ����   ����i�N  ����N  ���� +  ) g�1  i�N  ����N  ����i�   ����N  ����i�   ����   ����i�N  ����N  ���� /  ? g�1  i�N  ����N  ����i�   ����N  ����i�   ����   ����i�N  ����N  ���� 0  5 g�1  i�  4���N  4���i�  4���  4���i�N  4���N  4��� 8  C g�1  i��  4����  h���i��  4����  4���i�:  }���:  h���i�N  }���N  }���i��  h���:  h���i�:  }���N  }���i��  4����  4��� ,  4  : g�0 
 i��  �����  ����i��  T����  ����i��  �����  ����i�8  T����  T���i�N  ?���N  ?���i�8  ?���8  T���i��  �����  ����i��  �����  ����i��  �����  ����i�N  ?���8  ?��� 7 _   - g�1     $ 9  S g�1  i�  }����   }���i��   j����   }���i�  }���  }���i��   j���r  j���i�r  3���r  j���i�W  3���W  3���i�r  3���W  3���  =  % g�0  i��  �����  ����i��  �����  ����i��  �����  ����i��  �����  ���� [  1 g�0  i�a   f���a   f���i�a   f���Q   f���i�Q   f���Q   f��� d   3 < A  F g�0  i�d   ���d   ���i�d   ���S   ���i�S   ���S   ��� f  '  U g�Z       g�1  i��   ����  ����i��   �����   ����i�  ����  ����      Unknown Name