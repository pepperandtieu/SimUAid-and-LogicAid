�d d       d   " ��  Cclock   ����R   ����)   ����M   ����
 Clk       ��  CpinR   ����D   ����1 1 ClkR   ����        ��  CRegisterAdder%   ����m  G���                       �@   G���@   V���1 1 Clk6   G���        �X   ����X   ����0 0             LS    �?   ����?   ����0 0 Sh8   ����   RS    �m  q���^  q���0 0             Rin    �q   G���q   V���0 0                 ��   G����   V���1 1                 ��   G����   V���1 1                 �  G���  V���0 0                 �9  G���9  V���1 1                 �%   q���3   q���0 0 Add   ���   Ld    �%   d���3   d���0 0 LdM   q���   CLR    �Y   G���Y   V���0 0                   �Q  G���Q  V���0 0 P4B  G���        �   G���   V���0 0 P5  G���        ��   G����   V���0 0 P6�   G���        ��   G����   V���0 0 P7�   G���        ��   G����   V���0 0 P8�   G���                    nd   Register
for
Adder,  ����H  ����	   
                     ��  CShiftRegRS�  ����7  M���                      	 �  M���  [���1 1 Clk
  M���        ��  r����  r���0 0             Lin    ��  M����  [���1 1                 ��  M����  [���0 0                 ��  M����  [���1 1                 ��  M����  [���1 1                 �7  ~���)  ~���0 0 LdM:  ����   Ld    �7  r���)  r���0 0 Sh;  ~���   RS    �7  g���)  g���0 0             CLR     ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����0 0                              E(   Right
SRw   �����   ����            ����      �� 
 CNBitAdder�   :���m  ����                      	 �m  ���^  ���0 0             Cin    ��   :����   ,���0 0                 ��   :����   ,���0 0                 �   :���   ,���0 0                 �Q  :���Q  ,���0 0                 ��   �����   ����1 1                 ��   �����   ����1 1                 �  ����  ����0 0                 �F  ����F  ����1 1                  ��   :����   ,���1 1                  ��   :����   ,���1 1                  �  :���  ,���0 0                  �9  :���9  ,���1 1                  ��   ����   ���0 0             Cout                Ad   Adder
for
Register�   �����   ����������������          ��  Cswitch�   �����   �����   �����   ���� Mc1    ��   �����   ����1 ��                 ��   �����   ����0 ��                  ��   �����   ����1 1 Mc1�   ����        7��   �����   �����   �����   ���� Mc2    ��   �����   ����1 ��                 ��   �����   ����0 ��                  ��   �����   ����1 1 Mc2�   ����        7�  ����  ����  ����,  ���� Mc3    �  ����  ����1 ��                 �  ����  ����0 ��                  �  ����  ����0 0 Mc3  ����        7�>  ����J  ����5  ����_  ���� Mc4    �?  ����?  ����1 ��                 �K  ����K  ����0 ��                  �F  ����F  ����1 1 Mc45  ����        7��  K����  ����  ����  	��� Mp1    ��  ����  *���1 ��                 ��  ����  *���0 ��                  ��  M����  >���1 1 Mp1�  ���        7��  K����  ����  ����  	��� Mp2    ��  ����  *���1 ��                 ��  ����  *���0 ��                  ��  M����  >���0 0 Mp2�  ���        7��  K����  ����  ���  	��� Mp3    ��  ����  *���1 ��                 ��  ����  *���0 ��                  ��  M����  >���1 1 Mp3�  ���        7��  K���  ����  ���(  	��� Mp4    ��  ����  *���1 ��                 �  ���  *���0 ��                  ��  M����  >���1 1 Mp4�  ���        ��  Cground-  g���B  O���                          �7  g���7  X���0 0                  X�b  q���v  X���                          �m  q���m  c���0 0                  X�O   G���c   0���                          �Y   G���Y   :���0 0                  X�b   ����v   ����                          �l   ����l   ����0 0                  X�b  ���v  ����                          �m  ���m  ���0 0                  ��  CLoadableCounter�   �����   ����                       ��   �����   ����1 1 Clk�   ����        ��   �����   ����0 0 Sh�   ����   En    ��   �����   ����1 1             CLR     ��   �����   ����0 0                  ��   �����   ����0 0                  ��   �����   ����0 0              K                  (   CounterP   ����^   ����            �� 	 Cinverter�   ����2  ����                      �2  ����$  ����0 0                   ��   ����  ����1 1                  7�:   ���i   ���                       �:   ���G   ���1 ��                 �:   ���G   ���0 ��                  �i   	���\   	���0 0                  ��  CStateMachine�   i���  ���                       ��   ����   +���1 1 Clk�   ���        ��   ����   +���0 0 St�   ���       ��   ����   +���0 0 M�   ���       ��   ����   +���0 0 K�   ���        ��   i����   [���0 0 Sh�   v���        ��   i����   [���0 0 Add�   v���        ��   i����   [���0 0 Done�   ���        ��   i����   [���0 0 LdM�   w���                     E (   State
Machinew   �����   ������������               S0St'0S0S0StLdMS1S1K'M'ShS1S1K M'ShS3S1MAddS2S2K'ShS1S2KShS3S3-DoneS0��  CprobeH   ����\   ����U   ����y   ����  Clk     �R   ����R   ����1 1 ClkU   ����          }�f   >���z   ���Q   +���n   ���  St     �p   ���p   -���0 0 StQ   +���          }��   �����   �����   �����   ����  P8     ��   �����   ����0 0 P8�   ����          }��   �����   �����   �����   ����  P7     ��   �����   ����0 0 P7�   ����          }��   �����   �����   ����  ����  P6     ��   �����   ����0 0 P6�   ����          }�  ����*  ����$  ����E  ����  P5     �   ����   ����0 0 P5$  ����          }�F  ����Y  ����S  ����t  ����  P4     �O  ����O  ����0 0 P4S  ����          }��  �����  �����  �����  ����  P3     ��  �����  ����0 0 P3�  ����          }��  �����  �����  �����  ����  P2     ��  �����  ����0 0 P2�  ����          }��  �����  �����  ����  ����  P1     ��  �����  ����0 0 P1�  ����          }�  ����  ����
  ����%  ����  M     �  ����  ����0 0 M
  ����          }��   ����   �����   ����   ����  K     ��   �����   ���0 0 K�   ���          }��   �����   v����   �����   ����  Done     ��   v����   ����0 0 Done�   ����          & ��  Cnet1  ��  CsegmentR   ����R   ������R   ����R   ����    e u   ��1  ���   :����   G������   :����   :������   G����   G���   2 ��1  ���   :����   G������   :����   :������   G����   G���   3 ��0  ��  :���  G�����  :���  :�����  G���  G���   4 ��1  ��9  :���9  G�����9  :���9  :�����9  G���9  G���   5 ��1  ���   �����   �������   �����   ���� .  ; ��1  ���   �����   �������   �����   ���� /  ? ��0  ��  ����  ������  ����  ���� 0  C ��1  ��F  ����F  ������F  ����F  ���� 1  G ��1  ���  M����  M������  M����  M������  M����  M���   K ��0  ���  M����  M������  M����  M������  M����  M���   O ��1  ���  M����  M������  M����  M���   S ��1  ���  M����  M������  M����  M������  M����  M���   W ��0    	 ! f  y ��0  ��7  g���7  g�����7  g���7  g��� "  Z ��0  ��m  q���m  q�����m  q���m  q��� 
  \ ��0  ��Y   G���Y   G�����Y   G���Y   G���   ^ ��0  ��l   ����X   ������X   ����X   ������X   ����X   ������l   ����l   ����   ` ��0  ��m  ���m  �����m  ���m  ��� )  b ��0  ��q   G���q   ������   ���q   ������   ����   �����q   G���q   G���   6 ��0      z ��1  ���   �����   �������   �����   �������   �����   ���� g  n ��0  ���  �����  �������  �����  �������  �����  �������  �����  ���� �  # ��0  ���  �����  �������  �����  �������  �����  �������  �����  �������  �����  ���� �  $ ��0  ���  �����  �������  �����  �������  �����  �������  �����  �������  �����  ���� �  % ��0    �   ��0       ��0  ���   :����   :������   :����   G������   G����   G��� * �   ��0  ���   :����   :������   :����   G������   G����   G��� + �   ��0  ��   :���   :�����   :���   G�����   G���   G��� , �   ��0  ��Q  :���Q  :�����Q  :���Q  B�����Q  B���Q  G�����Q  B����  B������  r����  B������  r����  r������  r����  r�����Q  G���Q  G��� -  �   ��0  ���   i����   i������   i����   i������   v����   i������   v����   v������   v����   v��� �  { ��0  ���   	����   �����i   	���i   	������   ����   �����p   	����   	�����i   	���p   	�����p   	���p   �����p   ���p   ��� v �  r ��0  ��2  ����2  i������   i���2  i������   i����   i�����2  ����2  ���� m     | ��0  ���   �����   ������   �����   �������   ����   ������   �����   �������   �����   �������   �����   ���� x �  j ��X       ��0       ��0  ��  ����  ������  ����  �������  ����  �������  �����  ���� � w  &  ��  Ccomment
Multiplier�  ���  ����-�Multiplicand/   �����   ����-�Producth  �����  ����-�	(M is P0)  ����w  ����Tester using Debug version.