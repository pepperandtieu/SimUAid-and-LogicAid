�d d       d    ��  Cclock�   K���  :����   ]���  K���
 Clk       ��  Cpin  C���  C���1 1 Clk  Q���        ��  Cand3c   �����   ����                       �c   ����p   ����1 1 Sum2C   ����        �c   ����p   ����1 1 Sum1C   ����        �c   ����p   ����1 1 Sum0B   ����         ��   �����   ����1 1 D7�   ����        �a   �����   ����                       �a   ����p   ����0 0 Sum3A   ����        �a   ����p   ����1 1 Sum1A   ����        �a   ����p   ����1 1 Sum0A   ����         ��   �����   ����0 0                  ��  Cor2�   �����   ����                       ��   �����   ����1 1                  ��   �����   ����0 0                   ��   �����   ����1 1 D711�   ����        ��  Cxor20   c���s   >���                       �0   V���C   V���0 0 S3    `���        �0   J���C   J���0 0 Sum3   R���         �r   Q���d   Q���0 0                  �0   9���s   ���                       �0   .���C   .���0 0 S2    7���        �0   "���C   "���1 1 Sum2   *���         �r   (���d   (���1 1                  �0   ���s   ����                       �0    ���B    ���0 0 S1!   ���        �0   ����B   ����1 1 Sum1   ����         �r   ����d   ����1 1                  �/   ����r   ����                       �/   ����C   ����0 0 S0   ����        �/   ����C   ����1 1 Sum0   ����         �r   ����d   ����1 1                  �� 	 CbusinputQ  ^���m  A���^  |���v  j���  7       ��  Cbuspin^  ^���^  P���X X Sum@  e���         ��  �����  ����0 0 0�  ����        ��  �����  ����1 1 1�  ����        ��  �����  ����1 1 2�  ����        ��  �����  ����1 1 3�  ����                       �((       ����   ����            �� 	 Cinvertera   �����   k���                       �a   }���n   }���1 1 Sum2A   ����         ��   }����   }���0 0                  ��  Cnor4�   "����   ����                       ��   "����   "���0 0                  ��   ����   ���1 1                  ��   
����   
���1 1                  ��   �����   ����1 1                   ��   ����   ���0 0 Eq�   ���        ��   �����   q���                       ��   �����   ����0 0 Sum3�   ����        ��   }����   }���0 0                   ��   �����   ����0 0 D2312  ����        �� 	 CRegister  5����  ����                       �[  ����[  ����1 1 ClkQ  ����        ��  ���x  ���0 0 Sp�  #���   Ld    ��  ���x  ���0 0             CLR    �  ����  ����0 0 Sum3�   ����       �  ����  ����1 1 Sum2  ����       �2  ����2  ����1 1 Sum1$  ����       �E  ����E  ����1 1 Sum05  ����        �  5���  &���0 0 S3  B���        �  5���  &���0 0 S2  B���        �2  5���2  &���0 0 S1+  B���        �E  5���E  &���0 0 S0>  B���                     E (   Registerw   �����   ����         ��  CStateMachine#   �����   ?���                       ��   ?����   M���1 1 Clk�   ?���        �-   ?���-   M���0 0 Rb   B���       �@   ?���@   M���0 0 Reset/   A���       �T   ?���T   M���1 1 D7R   A���       �f   ?���f   M���1 1 D711Z   3���       �z   ?���z   M���0 0 D2312i   ?���       ��   ?����   M���0 0 Eq�   4���        �-   ����-   |���0 0 Sp!   ����        �@   ����@   |���0 0 Roll7   ����        �T   ����T   |���0 0 Win]   ����        �f   ����f   |���0 0 Loset   ����                      (   State
Machine�   �����   ����    ��n               S0Rb'0S0S0Rb0S1S1Rb' D7110S2S1RbRollS1S1Rb' D711' D23120S3S1Rb' D711' D2312'SpS4S2Reset'WinS2S2ResetWinS0S3Reset'LoseS3S3ResetLoseS0S4Rb'0S4S4Rb0S5S5Rb' Eq' D7'0S4S5RbRollS5S5
Rb' Eq' D70S3S5Rb' Eq0S2��  Cprobe�   �����   �����   �����   ����  Win     ��   �����   ����0 0 Win�   ����          W��   �����   �����   �����   ����  Lose     ��   �����   ����0 0 Lose�   ����          �� 	 CSplitter7  �����  l���                        (�^  l���^  z���Z Z                  �  ����  ����0 0 0�  ����        �  ����  ����1 1 1�  ����        �  ����  ����1 1 2�  ����        �  ����  ����1 1 3�  ����         �@  ����@  |���0 0 Sum30  ����        �T  ����T  |���1 1 Sum2F  ����        �h  ����h  |���1 1 Sum1Z  ����        �{  ����{  |���1 1 Sum0n  ����                      P(    O   ����O   ����O           ��  Cswitch'   0���3   ���!    ���C   ���� Rb    �'   ���'   ���1 Z                  �3   ���3   ���0 Z                   �-   0���-   #���0 0 Rb!    ���        g�C   .���P   ����A   ����v   ���� Reset    �C   ����C   ���1                    �P   ����P   ���0 1                   �I   .���I   !���0 0 ResetA   ����        ��  Cground�  ����  ����                          ��  ����  ����0 0                   ��  CbusZ       ��  Cnet0  ��  Csegment�   �����   ����w��   �����   ����w��   �����   ����w��   �����   ����    u�1  w��   �����   ����w��   �����   ����w��   �����   ����w��   �����   ����  O  
 u�1  w�r   ����r   ����w��   
����   
���w�r   
����   
���w�r   ����r   
��� 6  ! u�1  w�r   (���r   (���w��   ����   ���w�r   ����   ���w�r   (���r   ��� 5   s�Z       u�0  w��   }����   }���w��   }����   }���w��   }����   }��� ;  1 u�1      0 C  d u�1        D  e u�1  w��   �����   ����w�r   ����r   ����w��   �����   ����w�r   �����   ���� 7  % u�0  w�r   Q���r   Q���w��   "����   "���w�r   Q����   Q���w��   "����   Q��� 4   u�1    	  $ E  f u�0      : B  c u�1    P   u�0  w��  ����  ���w��  ����  ���w��  ����  ���w��  ����  ��� A  r u�0  w�T   ����T   ����w�T   ����T   ����w�T   �����   ����w��   �����   ����w��   �����   ���� Y  U u�0  w��   �����   ����w�f   �����   ����w�f   ����f   ����w��   �����   ���� [  V u�0      F u�Z  w��  �����  ����    s�Z  w�^  l���^  l���w�^  ^���^  ^���w�^  ^���^  l��� ^  ) u�0  w�-   0���-   0���w�-   ?���-   ?���w�-   0���-   ?��� M  k u�0  w�@   2���@   ?���w�@   ?���@   ?���w�I   .���I   .���w�I   2���I   .���w�I   2���@   2��� N  o u�0      G u�0      H u�0    #  I u�0    R  8 u�0    Q  < u�0    @  S u�0       u�0       u�1    ? L     Dr. Charles Roth      