�d d        d    ��  CRegisterAdder�   a����  ���                       ��  Cpin�   ����   ���0 0 Clk�   ���        ��   a����   S���0 0             LS    ��   a����   S���0 0 Sh�   m���   RS    ��  8����  8���0 0             Rin    ��   ����   ���0 0                 �!  ���!  ���0 0                 �S  ���S  ���0 0                 ��  ����  ���0 0                 ��  ����  ���0 0                 ��   9����   9���0 0 Add�   E���   Ld    ��   ,����   ,���0 0 LdM�   8���   CLR    ��   ����   ���0 0                   ��  ����  ���0 0 P4�  ���        ��  ����  ���0 0 P5�  ���        �l  ���l  ���0 0 P6e  ���        �:  ���:  ���0 0 P73  ���        �  ���  ���0 0 P8  ���                    nd   Register
for
Adder,  ����H  ����	   
                     �� 
 CNBitAdder  ����  ����                      	 ��  �����  ����0 0             Cin    �:  ���:  ����0 0                 �l  ���l  ����0 0                 ��  ����  ����0 0                 ��  ����  ����0 0                 �.  ����.  ����0 0                 �`  ����`  ����0 0                 ��  �����  ����0 0                 ��  �����  ����0 0                  �!  ���!  ����0 0                  �S  ���S  ����0 0                  ��  ����  ����0 0                  ��  ����  ����0 0                  �  ����  ����0 0             Cout                Ad   Adder
for
Register�   �����   ���� 3   h/           ��  Cground�  8����   ���                          ��  8����  *���0 0                  %��   ����   ����                          ��   ����   ����0 0                  %��   m���  U���                          ��   m����   _���0 0                  %��  �����  ����                          ��  �����  ����0 0                  ��  CShiftRegRS  W����  ���                      	 ��  ����  ���0 0 Clk�  ���        �  1���(  1���0 0             Lin    �2  ���2  ���0 0                 �F  ���F  ���0 0                 �Z  ���Z  ���0 0                 �n  ���n  ���0 0                 ��  =����  =���0 0 LdM�  I���   Ld    ��  1����  1���0 0 Sh�  =���   RS    ��  %����  %���0 0             CLR     �2  W���2  I���0 0 P3+  d���        �F  W���F  I���0 0 P2?  d���        �Z  W���Z  I���0 0 P1S  d���        �n  W���n  I���0 0 Mk  e���                    E(   Right
SRx   �����   ����            ����      %��  %����  ���                          ��  %����  ���0 0                  ��  Cprobe�   ����  �����   ����  ����  P8     ��   �����   ����0 0 P8�   ����          ?�  ����,  ����  ����:  ����  P7     �"  ����"  ����0 0 P7  ����          ?�>  ����R  ����?  ����`  ����  P6     �H  ����H  ����0 0 P6?  ����          ?�c  ����w  ����a  �����  ����  P5     �m  ����m  ����0 0 P5a  ����          ?��  �����  �����  �����  ����  P4     ��  �����  ����0 0 P4�  ����          ?��  �����  �����  �����  ����  P3     ��  �����  ����0 0 P3�  ����          ?��  �����  �����  �����  ����  P2     ��  �����  ����0 0 P2�  ����          ?�  ����  ����  ����'  ����  P1     �  ����  ����0 0 P1  ����          ?�/  ����C  ����2  ����K  ����  M     �9  ����9  ����0 0 M2  ����          ��  CswitchZ   �����   ����g   �����   ���� Sh     �Z   ����h   ����1                    �Z   ����h   ����0 '                   ��   ����|   ����0 0 Shg   ����        R�V   �����   ����c   �����   ���� Add     �V   ����d   ����1                    �V   ����d   ����0                     ��   ����x   ����0 0 Addc   ����        R�U   Y����   M���_   r����   `��� Clk     �U   Y���c   Y���1                   �U   M���c   M���0                    ��   S���w   S���0 0 Clk_   r���        R��   ����.  ����  ����4  ���� Mc3     ��   ����  ����1                    ��   ����  ����0                     �.  ����   ����0 0 Mc3  ����        R�0  }���`  q���=  ����f  }��� Mc2     �0  }���>  }���1 ��                 �0  q���>  q���0 1                   �`  w���R  w���0 0 Mc2=  ����        R�T  [����  O���a  m����  [��� Mc1     �T  [���b  [���1                    �T  O���b  O���0                     ��  U���v  U���0 0 Mc1a  m���        R��  ;����  /����  M����  ;��� Mc0     ��  ;����  ;���1 ��                 ��  /����  /���0                     ��  5����  5���0 0 Mc0�  M���        R�  ����3  ����  
���9  ���� Mp3     �  ����  ����1 ��                 �  ����  ����0                    �3  ����%  ����0 0 Mp3  
���        R�  ����G  ����$  ����M  ���� Mp2     �  ����%  ����1                    �  ����%  ����0 ��                  �G  ����9  ����0 0 Mp2$  ����        R�*  ����Z  ����7  ����`  ���� Mp1     �*  ����8  ����1                    �*  ����8  ����0 ��                  �Z  ����L  ����0 0 Mp17  ����        R�>  ����n  ����K  ����t  ���� Mp0     �>  ����L  ����1                    �>  ����L  ����0                     �n  ����`  ����0 0 Mp0K  ����        R�Y   �����   |���f   �����   ���� LdM     �Y   ����g   ����1                    �Y   |���g   |���0 ��                  ��   ����{   ����0 0 LdMf   ����          ��  Cnet0  ��  Csegment!  ���!  �����!  ���!  �����!  ���!  ��� 	    ��0  ��S  ���S  �����S  ���S  �����S  ���S  ��� 
  ! ��0  ���  ����  ������  ����  ������  ����  ���   " ��0  ���  ����  ������  ����  ������  ����  ���   # ��0  ���   ����   �����  ����  �������   �����   �����  �����   ����   $ ��0  ���  8����  8������  8����  8������  8����  8���   ' ��0  ���   ����   ������   ����   ������   ����   ���   ) ��0  ���  �����  �������  �����  �������  �����  ����   - ��0     0  ^ ��0  ���   a����   a������   m����   m������   m����   a������   m����   m���   + ��0  ���  %����  %������  %����  %������  %����  %��� 8  > ��0     7  V ��0      Z ��0     6  � ��0    A   ��0  ��:  ���:  �����:  ���:  �����:  ���:  ���  C   ��0  ��l  ���l  �����l  ���l  �����l  ���l  ���  E   ��0  ���  ����  ������  ����  ������  ����  ���  G   ��0  ���  ����  ������  ����  �����  ����  �����  1���  1������  ����  �����  1���  ���  1 I   ��0    K  9 ��0    M  : ��0    O  ; ��0    Q  < ��0  ��.  ����.  ������.  ����.  ������.  ����.  ����   b ��0  ��`  ����`  ������`  w���`  w�����`  w���`  ����   f ��0  ���  �����  �������  U����  U������  U����  �������  U����  U���   j ��0  ���  �����  �������  5����  5������  5����  �������  5����  5���   n ��0  ��2  ���2  �����3  ����3  ������3  ���2  �����3  ����3  ��� 2  r ��0  ��F  ���F  �����G  ����G  ������F  ����F  �����G  ����F  ���� 3  v ��0  ��Z  ���Z  �����Z  ����Z  ������Z  ����Z  ��� 4  z ��0  ��n  ���n  �����n  ����n  ������n  ����n  ��� 5  ~ ��0        ��  CcommentMultiplicandA  $����  �����
Multiplier&  �����  i���Dr. Charles Roth      