 �d d       d    ��  Cclock�   \����   J����   n����   \���
 clock       ��  Cpin�   T����   T���0 1 clock�   b���        ��  CBShiftRegLS�   ����x  h���                       �  h���  v���0 0                  �x  ����j  ����0 0             Rin    ��  CbuspinC  h���C  v���Z Z                 	 �w  4���w  B���1 1 0t  4���        �w  4���w  B���1 1 1t  4���        �w  4���w  B���0 0 2t  4���        �w  4���w  B���0 0 3t  4���        �w  4���w  B���0 0 4t  4���        �w  4���w  B���1 1 5t  4���        �w  4���w  B���0 0 6t  4���        �w  4���w  B���1 1 7t  4���        �w  4���w  B���1 1 8t  4���        ��   �����   ����0 0             Ld    ��   �����   ����0 0 Sh�   ����   LS    ��   �����   ����0 0             CLR     	�C  ����C  ����X X                  	 �w  ����w  r���0 0 0t  ����        �w  ����w  r���0 0 1t  ����        �w  ����w  r���1 1 2t  ����        �w  ����w  r���0 0 3t  ����        �w  ����w  r���1 1 4t  ����        �w  ����w  r���1 1 5t  ����        �w  ����w  r���0 0 6t  ����        �w  ����w  r���1 1 7t  ����        �w  ����w  r���0 0 8t  ����                    	F!(   Left
SRv   �����   ����                ����   �� 
 CBNWideMux�   Z����  ���                       �  5���  5���0 0 Load�   =���   S    	�/  ���/  ���Z Z                 	 �c  ����c  ����1 1 0`  ����        �c  ����c  ����1 1 1`  ����        �c  ����c  ����0 0 2`  ����        �c  ����c  ����0 0 3`  ����        �c  ����c  ����0 0 4`  ����        �c  ����c  ����1 1 5`  ����        �c  ����c  ����0 0 6`  ����        �c  ����c  ����1 1 7`  ����        �c  ����c  ����1 1 8`  ����        	�W  ���W  ���Z Z                 	 ��  �����  ����0 0 0�  ����        ��  �����  ����1 1 1�  ����        ��  �����  ����0 0 2�  ����        ��  �����  ����0 0 3�  ����        ��  �����  ����0 0 4�  ����        ��  �����  ����0 0 5�  ����        ��  �����  ����1 1 6�  ����        ��  �����  ����1 1 7�  ����        ��  �����  ����1 1 8�  ����         	�C  Z���C  L���X X                  	 �w  ���w  ����1 1 0t  ���        �w  ���w  ����1 1 1t  ���        �w  ���w  ����0 0 2t  ���        �w  ���w  ����0 0 3t  ���        �w  ���w  ����0 0 4t  ���        �w  ���w  ����1 1 5t  ���        �w  ���w  ����0 0 6t  ���        �w  ���w  ����1 1 7t  ���        �w  ���w  ����1 1 8t  ���                    	!(   
2-to-1
Muxw   �����   ����         �� 
 CBusMergerh  �����  ����                        	�r  ����r  ����Z Z             1    ��  �����  ����0 0                  	��  �����  ����Z Z             8    ��  �����  ����1 1                  ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                   	�|  ����|  ����X X             9    	 ��  �����  ����0 0                  ��  �����  ����1 1                  ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                                	�(    (   ����(   ��������   ������  CComplementer�   M���  ���                       ��   '����   '���1 1                  	��   ����   ���Z Z                  �	  v���	  ����0 0 0  v���        �	  v���	  ����1 1 1  v���        �	  v���	  ����1 1 2  v���        �	  v���	  ����0 0 3  v���        �	  v���	  ����1 1 4  v���         	��   M����   ?���X X                   �	  ����	  ����1 1 0  ����        �	  ����	  ����0 0 1  ����        �	  ����	  ����0 0 2  ����        �	  ����	  ����1 1 3  ����        �	  ����	  ����0 0 4  ����                    B`(   Complementerc   ����   ����O           B��   ����4  ����                        	�  ����  ����Z Z             5    �6  i���6  w���1 1                  �6  i���6  w���1 1                  �6  i���6  w���0 0                  �6  i���6  w���0 0                  �6  i���6  w���0 0                  	�  ����  ����Z Z             3    �J  ����J  ����1 1                  �J  ����J  ����0 0                  �J  ����J  ����1 1                  	�*  ����*  ����Z Z             1    �*  ����*  ����1 1                   	�  ����  ����X X             9    	 �J  ����J  ����1 1                  �J  ����J  ����1 1                  �J  ����J  ����0 0                  �J  ����J  ����0 0                  �J  ����J  ����0 0                  �J  ����J  ����1 1                  �J  ����J  ����0 0                  �J  ����J  ����1 1                  �J  ����J  ����1 1                                	�(    ;   ����;   ���� CLR     B��   �����   ����                        	��   �����   ����Z Z             1    �   ����   ����0 0                  	��   �����   ����Z Z             4    �  ����  ����1 1                  �  ����  ����1 1                  �  ����  ����0 0                  �  ����  ����1 1                   	��   �����   ����X X             5     �
  ����
  ~���0 0                  �
  ����
  ~���1 1                  �
  ����
  ~���1 1                  �
  ����
  ~���0 0                  �
  ����
  ~���1 1                                �(    (   ����(   �����6  i���6��  CBusSplitter�   y���4  I���                        	�  I���  W���Z Z                 	 �U  9���U  G���0 0 0R  9���        �U  9���U  G���0 0 1R  9���        �U  9���U  G���1 1 2R  9���        �U  9���U  G���0 0 3R  9���        �U  9���U  G���1 1 4R  9���        �U  9���U  G���1 1 5R  9���        �U  9���U  G���0 0 6R  9���        �U  9���U  G���1 1 7R  9���        �U  9���U  G���0 0 8R  9���         	�  y���  k���X X             5     �A  j���A  \���0 0                  �A  j���A  \���0 0                  �A  j���A  \���1 1                  �A  j���A  \���0 0                  �A  j���A  \���1 1                  	�  y���  k���X X             3     �U  j���U  \���1 1                  �U  j���U  \���0 0                  �U  j���U  \���1 1                  	�*  y���*  k���X X X0#  ����   1     �i  j���i  \���0 0                                	�(    ;   ����;   �������   �  ��  Cgroundh  ����|  ����                          �r  ����r  ����0 0                  ���   �����   ����                          ��   �����   ����0 0                  ��  CplusVB  ����V  ����                          �K  ����K  ����1 1                  �� 	 Cbusinputt  �����  �����  �����  ����  87       	��  �����  ����X X dividendl  ����         ��  �����  ����1 1 0�  ����        ��  �����  ����0 0 1�  ����        ��  �����  ����0 0 2�  ����        ��  �����  ����0 0 3�  ����        ��  �����  ����0 0 4�  ����        ��  �����  ����1 1 5�  ����        ��  �����  ����1 1 6�  ����        ��  �����  ����1 1 7�  ����                       �((    $   ����$   �����           ���   �����   �����   7���  %���  d       	��   �����   ����X X divisor�   ����         �  ����  ����1 1 0  ����        �  ����  ����1 1 1  ����        �  ����  ����0 0 2  ����        �  ����  ����1 1 3  ����                       �((       ����   �����           ��  Cor2�   �����   ����                       ��   �����   ����0 0 Loadi   ����        ��   �����   ����0 0 Suv   ����         ��   �����   ����0 0                  ��}  �����  l���                          ��  �����  v���0 0                  ��R  �����  \���                        	�p  \���p  j���Z Z                 	 �v  Z���v  h���0 0 0s  Z���        �v  Z���v  h���0 0 1s  Z���        �v  Z���v  h���1 1 2s  Z���        �v  Z���v  h���0 0 3s  Z���        �v  Z���v  h���1 1 4s  Z���        �v  Z���v  h���1 1 5s  Z���        �v  Z���v  h���0 0 6s  Z���        �v  Z���v  h���1 1 7s  Z���        �v  Z���v  h���0 0 8s  Z���         	�\  ����\  ~���X X             1     �b  ����b  }���0 0                  	�p  ����p  ~���X X             4     �v  ����v  }���0 0                  �v  ����v  }���1 1                  �v  ����v  }���0 0                  �v  ����v  }���1 1                  	��  �����  ~���X X             4     ��  �����  }���1 1                  ��  �����  }���0 0                  ��  �����  }���1 1                  ��  �����  }���0 0                                	�(    ;   ����;   ����        6   �� 	 Cbusprobe.  ����I  ����  ����m  ����  	remainder     	�<  ����<  ����Z Z 	remainder  ����         �^  ����^  ����0 0 0[  ����        �^  ����^  ����1 1 1[  ����        �^  ����^  ����0 0 2[  ����        �^  ����^  ����1 1 3[  ����                          H(       ����   �������{   n  ܀�  �����  �����  �����  ����  quotient     	��  �����  ����Z Z quotient�  ����         ��  �����  ����1 1 0�  ����        ��  �����  ����0 0 1�  ����        ��  �����  ����1 1 2�  ����        ��  �����  ����0 0 3�  ����                          H(       ����   ����        ��  CStateMachineK   ,����   ����                       ��   �����   ����0 0 clock�   ����        �T   ����T   ����1 1 St?   ����       �h   ����h   ����0 0 Cm   ����        �T   ,���T   ���0 0 Load=   ;���        �h   ,���h   ���0 0 Sha   ;���        �|   ,���|   ���0 0 Suu   ;���        ��   ,����   ���0 0 V�   ;���                     E (   State
Machinev   �����   ������������               S0St'0S0S0StLoadS1S1CVS0S1C'ShS2S2CSuS2S2C'ShS3S3CSuS3S3C'ShS4S4CSuS4S4C'ShS5S5CSuS0S5C'0S0���   �����   h���                          ��   �����   r���0 0                  ��  CswitchM   ����Y   ����                      �O   ����O   ����1 ��                 �Z   ����Z   ����0 ��                  �T   ����T   ����1 1                  ��  CBNBitAdderCluster   ����  Y���                       �  ����   ���1 1             Cin    	��   Y����   g���Z Z                  ��   R����   `���0 0 0�   R���        ��   R����   `���0 0 1�   R���        ��   R����   `���1 1 2�   R���        ��   R����   `���0 0 3�   R���        ��   R����   `���1 1 4�   R���        	��   Y����   g���Z Z                  ��   R����   `���1 1 0�   R���        ��   R����   `���0 0 1�   R���        ��   R����   `���0 0 2�   R���        ��   R����   `���1 1 3�   R���        ��   R����   `���0 0 4�   R���         	��   �����   ����X X                   ��   �����   ����1 1 0�   ����        ��   �����   ����1 1 1�   ����        ��   �����   ����0 0 2�   ����        ��   �����   ����0 0 3�   ����        ��   �����   ����0 0 4�   ����        �   ����   ���0 0             Cout                A2   Adderp   ������/ ��/ ��/  �/ ��/            ��  CbusZ  ��  CsegmentC  Z���C  h����C  Z���C  Z����C  h���C  h��� 
  8 �Z  �W  ����W  ����|  ����|  �����W  ���W  ����|  ����|  �����|  ����W  ���� .  O �Z  ��   M����   M�����   Y����   Y�����   Y����   M���  b �Z  �/  ���/  ����  ����  �����/  ���/  ����  ����  ����  ���/  ��� $  u �Z  �  ����  �����  ����  ������   ����  ������   �����   ������   �����   ���� i  �Z  ��   �����   ������   ����   �����   �����   ��� \  � �Z  �  y���  y����{   y���{   L�����   L���{   L����  y���{   y�����   Y����   Y�����   Y����   L��� �  � �Z  �  y���  �����  y���  y����  ����  ���� o  � �Z  �C  ����C  �����  ����C  �����C  ����C  �����  9���  �����  I���  D����  I���  I����  D���  D����  D���  9����  9���p  9����p  \���p  9����p  \���p  \��� � �   ��  Cnet0  �r  ����r  �����r  ����r  �����r  ����r  �����r  ����r  ���� D  � F�0  ��   �����   ������   �����   ������   �����   ������   �����   ���� �  � �Z  ��  �����  ������  �����  ������  �����  ���� F  � �Z  ��   �����   ������   �����   ������   �����   ���� �  � F�0  ��   �����   ������   �����   ������   �����   ������   �����   ����   � F�0  ��  �����  �����x  �����  �����x  ����x  ������  �����  ����   � F�0      � �Z  ��  �����  ������  �����  ������  �����  ������  �����  ������  �����  ���� �  � �Z  �p  ����p  �����<  ����<  �����p  ����p  �����<  ����p  �����<  ����<  ���� �  � F�0  ��   �����   ������   �����   ������   �����   ����   � F�0    # �  � F�0    �  � F�1  �T   ����T   �����T   ����T   �����T   ����T   ���� �  � F�0  �  h���  h����  h���  T�����   T���  T�����   T����   T���  �   F�1  �  ���K  ����K  ����K  ����K  ����K  �����  ���  ����K  ����K  �����K  ����*  �����*  ����*  �����*  ����*  ���� � s  � F�0  �   ���h   ����h   ����h   ����h   ����h   �����   ���   ��� �    testing               