 �d d         <    ��  Cclockn   �����   ����m   �����   ���� Clock       ��  Coutput�   �����   ����1 0 Clockm   ����        ��  CJKflipflop�   ����*  ^���                       ��  Cinput�   �����   ����1 1                  ��   �����   ����0 0                  ��   ~����   ~���1 1                  �  ����  ����1 1                  �  ^���  l���1 1                   �*  ����  ����0 0                  �*  ����  ����1 1                  ��   >���*  ����                       ��   ����   ���1 1                  ��   ����   ���1 1                  ��   �����   ����1 1                  �  >���  1���1 1                  �  ����  ����1 1                   �*  ���  ���0 0                  �*  ���  ���1 1                  ��  Cand2�   �����   ����                       ��   �����   ����0 0                  ��   �����   ����1 1                   ��   �����   ����0 0                  ��   1����   ���                       ��   %����   %���1 1                  ��   ����   ���1 1                   ��   ����   ���1 1                  ��  Cinput_signal   ����=   ����   ����.   ���� X       �=   ����/   ����1 1 X   ����         ��  Csignal    1 #�   0 #�    1 ��  Cxor2N  ����  ����                       �N   ���a   ���0 0                  �N  ����a  ����1 1                   ��  �����  ����1 1                  ��  Cswitch�   ����  �����   ����  ���� S1     ��   �����   ����1 Z                  ��   �����   ����0 Z                   �  �����   ����1 1 S1�   ����        ,��   ����'  ����  ����  ���� R     ��   ����  ����1 Z                  ��   ����  ����0 Z                   �'  ����  ����1 1 R  ����        ,��   C���	  7����   U���  C��� S2     ��   C����   C���1 Z                  ��   7����   7���0 Z                   �	  =����   =���1 1 S2�   U���        ��  Cprobe�   �����   �����   �����   ����  Clock     ��  Cpin�   �����   ����1 1 Clock�   ����          9�1   ����E   ����>   ����W   ����  X     ;�;   ����;   ����1 1 X>   ����          9�X  ����l  ����e  �����  ����  Q1     ;�b  ����b  ����0 0 Q1e  ����          9�N  F���b  &���[  X���|  F���  Q2     ;�X  &���X  4���0 0 Q2[  X���          9��  !����  ����  3����  !���  Z     ;��  ����  ���1 1 Z�  3���           ��  Cnet0  ��  Csegment�   �����   ����G��   �����   ����G��   �����   ���� 	   E�1  G��   ����   ���G��   ����   ���G��   ����   ���    E�1  G�*  ����*  ����G�o   T���o   %���G��   %����   %���G�o   %����   %���G�*  T���o   T���G�*  ����*  T���    E�1  G�=   ����=   ����G��   �����   ����G�M   ~���M   ���G��   ���M   ���G��   ����   ���G�M   ����M   ~���G��   ~����   ~���G�M   ���M   ����G��   ����M   ����G��   �����   ����G�M   ����M   ����G�N  ����N  ����G�N  ����N  ����G�M   ����N  ����G��   ~���M   ~���G��   ����M   ����G�=   ����M   ����G�;   ����=   ����G�;   ����;   ����   
  * >  " E�Z       E�1 
 G��   �����   ����G��   �����   ���G��   �����   ����G��   ����   ���G��   �����   ���G��   ����   ���G��   �����   ����G��   �����   ����G��   �����   ����G��   �����   ����   <   E�1  G�  ����  ����G�  ����  ����G�  ����  ����G�  ����  ����   0 E�1 	 G�  ^���  ^���G�&  ����'  ����G�'  ����'  ����G�&  ����&  ����G�  ����  ����G�&  ����  ����G�3  ����&  ����G�3  ^���  ^���G�3  ����3  ^���    4 E�1  G�  >���	  >���G�	  =���	  >���G�	  =���	  =���G�  >���  >���   8 E�0  G��   �����   ����G��   �����   ����G�=  �����   ����G�=  ����=  ���G�=  ���*  ���G�X  ���=  ���G�=  ���=   ���G�N   ���=   ���G�N   ���N   ���G�*  ���*  ���G�X  &���X  &���G�X  &���X  ���  ) B   E�1  G��  ����  ���G��  �����  ����G��  �����  ����G��  ����  ���� D  + E�0  G�b  ����b  ����G�*  ����b  ����G�*  ����*  ����G�b  ����b  ���� @     Unknown Name