�l l        d    ��  CBShiftRegLS�   ����c  W���                       ��  Cpin�   W����   e���1 1 clock�   [���        �c  ���T  ���0 0             Rin    ��  Cbuspin*  W���*  e���Z Z                 	 �w  4���w  B���1 1 0t  4���        �w  4���w  B���0 0 1t  4���        �w  4���w  B���0 0 2t  4���        �w  4���w  B���0 0 3t  4���        �w  4���w  B���1 1 4t  4���        �w  4���w  B���0 0 5t  4���        �w  4���w  B���0 0 6t  4���        �w  4���w  B���0 0 7t  4���        �w  4���w  B���1 1 8t  4���        ��   �����   ����1 1             Ld    ��   ����   ���0 0             LS    ��   r����   r���0 0             CLR     �*  ����*  ����X X                  	 �w  ����w  r���0 0 0t  ����        �w  ����w  r���0 0 1t  ����        �w  ����w  r���0 0 2t  ����        �w  ����w  r���0 0 3t  ����        �w  ����w  r���0 0 4t  ����        �w  ����w  r���0 0 5t  ����        �w  ����w  r���0 0 6t  ����        �w  ����w  r���0 0 7t  ����        �w  ����w  r���0 0 8t  ����                    	F!+   Left
SR�   �����   ����                ����   �� 
 CBNWideMux�   H���y  ����                       ��    ����    ���0 0 Load�   (���   S    �  ����  ���Z Z                 	 �c  ����c  ����1 1 0`  ����        �c  ����c  ����0 0 1`  ����        �c  ����c  ����0 0 2`  ����        �c  ����c  ����0 0 3`  ����        �c  ����c  ����1 1 4`  ����        �c  ����c  ����0 0 5`  ����        �c  ����c  ����0 0 6`  ����        �c  ����c  ����0 0 7`  ����        �c  ����c  ����1 1 8`  ����        �?  ����?  ���Z Z                 	 ��  �����  ����0 0 0�  ����        ��  �����  ����1 1 1�  ����        ��  �����  ����1 1 2�  ����        ��  �����  ����0 0 3�  ����        ��  �����  ����1 1 4�  ����        ��  �����  ����1 1 5�  ����        ��  �����  ����1 1 6�  ����        ��  �����  ����1 1 7�  ����        ��  �����  ����1 1 8�  ����         �*  H���*  9���X X                  	 �w  ���w  ����1 1 0t  ���        �w  ���w  ����0 0 1t  ���        �w  ���w  ����0 0 2t  ���        �w  ���w  ����0 0 3t  ���        �w  ���w  ����1 1 4t  ���        �w  ���w  ����0 0 5t  ���        �w  ���w  ����0 0 6t  ���        �w  ���w  ����0 0 7t  ���        �w  ���w  ����1 1 8t  ���                    	!+   
2-to-1
Mux�   �����   ����         �� 
 CBusMergerR  ����}  ����                        �]  ����]  ����Z Z             1    ��  �����  ����0 0                  �r  ����r  ����Z Z             8    ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����0 0                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                   �g  ����g  ����X X             9    	 ��  �����  ����0 0                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����0 0                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                                	�+    +   ����+   ��������   ������  CBNBitAdderClusterW   �����   /���                       ��   X����   X���1 1             Cin    ��   /����   >���Z Z                  ��   �����   ����0 0 0�   ����        ��   �����   ����0 0 1�   ����        ��   �����   ����0 0 2�   ����        ��   �����   ����0 0 3�   ����        ��   �����   ����0 0 4�   ����        ��   /����   >���Z Z                  �
  ����
  ����1 1 0  ����        �
  ����
  ����0 0 1  ����        �
  ����
  ����0 0 2  ����        �
  ����
  ����0 0 3  ����        �
  ����
  ����0 0 4  ����         ��   �����   r���X X                   ��   3����   %���1 1 0�   ?���        ��   3����   %���0 0 1�   ?���        ��   3����   %���0 0 2�   ?���        ��   3����   %���0 0 3�   ?���        ��   3����   %���1 1 4�   ?���        �W   X���f   X���0 0             Cout                Al   Adderx   �����   ����                     ��  CComplementerq   %����   ����                       �q   �����   ����1 1                  ��   �����   ����Z Z                  �	  v���	  ����0 0 0  v���        �	  v���	  ����1 1 1  v���        �	  v���	  ����1 1 2  v���        �	  v���	  ����1 1 3  v���        �	  v���	  ����1 1 4  v���         ��   %����   ���X X                   �	  ����	  ����1 1 0  ����        �	  ����	  ����0 0 1  ����        �	  ����	  ����0 0 2  ����        �	  ����	  ����0 0 3  ����        �	  ����	  ����0 0 4  ����                    B`+   Complementerk   �����   ����O           ?��   ����  ����                        ��   �����   ����Z Z             5    �6  i���6  w���1 1                  �6  i���6  w���0 0                  �6  i���6  w���0 0                  �6  i���6  w���0 0                  �6  i���6  w���1 1                  ��   �����   ����Z Z             3    �J  ����J  ����0 0                  �J  ����J  ����0 0                  �J  ����J  ����0 0                  �  ����  ����Z Z             1    �X  ����X  ����1 1                   ��   �����   ����X X             9    	 �J  ����J  ����1 1                  �J  ����J  ����0 0                  �J  ����J  ����0 0                  �J  ����J  ����0 0                  �J  ����J  ����1 1                  �J  ����J  ����0 0                  �J  ����J  ����0 0                  �J  ����J  ����0 0                  �J  ����J  ����1 1                                	�+    @   ����@   ���� CLR     ?��   �����   ����                        ��   �����   ����Z Z             1    �   ����   ����0 0                  ��   �����   ����Z Z             4    �  ����  ����1 1                  �  ����  ����1 1                  �  ����  ����1 1                  �  ����  ����1 1                   ��   �����   ����X X             5     �
  ����
  ~���0 0                  �
  ����
  ~���1 1                  �
  ����
  ~���1 1                  �
  ����
  ~���1 1                  �
  ����
  ~���1 1                                �+    +   ����+   �����6  i���6��  CBusSplitter�   @���  ���                        ��   ����   ���Z Z                 	 �U  9���U  G���0 0 0R  9���        �U  9���U  G���0 0 1R  9���        �U  9���U  G���0 0 2R  9���        �U  9���U  G���0 0 3R  9���        �U  9���U  G���0 0 4R  9���        �U  9���U  G���0 0 5R  9���        �U  9���U  G���0 0 6R  9���        �U  9���U  G���0 0 7R  9���        �U  9���U  G���0 0 8R  9���         ��   @����   1���X X             5     �A  j���A  \���0 0                  �A  j���A  \���0 0                  �A  j���A  \���0 0                  �A  j���A  \���0 0                  �A  j���A  \���0 0                  ��   @����   1���X X             3     �U  j���U  \���0 0                  �U  j���U  \���0 0                  �U  j���U  \���0 0                  �  @���  1���X X X0  S���   1     �i  j���i  \���0 0                                	�+    A   ����A   �������   �  ��  CgroundR  ����g  t���                          �]  ����]  ���0 0                  ���   �����   s���                          ��   �����   ~���0 0                  ��  CplusV)  ����>  ����                          �2  ����2  ����1 1                  �� 	 Cbusinput_  x����  W���m  �����  ����  DF       �r  x���r  i���X X dividendY  S���         ��  �����  ����1 1 0�  ����        ��  �����  ����1 1 1�  ����        ��  �����  ����0 0 2�  ����        ��  �����  ����1 1 3�  ����        ��  �����  ����1 1 4�  ����        ��  �����  ����1 1 5�  ����        ��  �����  ����1 1 6�  ����        ��  �����  ����1 1 7�  ����                       �(+    '   ����'   �����           ���   {����   Y����   ����   ����  F       ��   {����   k���X X divisor�   W���         �  ����  ����1 1 0  ����        �  ����  ����1 1 1  ����        �  ����  ����1 1 2  ����        �  ����  ����1 1 3  ����                       �(+       ����   �����           ��  Cor2a   �����   ����                       �a   ����u   ����0 0                  �a   ����u   ����1 1                   ��   �����   ����1 1                  ��  Cswitch   ����H   ����!   ����W   ���� Load     �   ����$   ����1 X                  �   ����$   ����0 Z                   �H   ����9   ����0 0 Load!   ����        ր   ����G   ����"   ����G   ���� Su     �   ����"   ����1                   �   ����"   ����0                     �G   ����8   ����1 1 Su"   ����        ր   ����G   y���"   ����G   ���� Sh     �   ����"   ����1                    �   y���"   y���0                    �G   ����8   ����0 0 Sh"   ����        ր   Y���G   L���"   l���H   Y��� Clr     �   Y���"   Y���1                    �   L���"   L���0                     �G   S���8   S���0 0 Clr"   l���        ր   -���H    ���"   C���X   0��� clock     �   -���$   -���1 z                  �    ���$    ���0 z                   �H   &���9   &���1 1 clock"   C���        ��h  u���~  [���                          �s  u���s  f���0 0                  ��  Cprobe   ����$   }���   ����P   ����  carry     �   }���   ����0 0 carry   ����          ��O  ~����  J���                        �o  J���o  Y���Z Z                 	 �v  Z���v  h���0 0 0s  Z���        �v  Z���v  h���0 0 1s  Z���        �v  Z���v  h���0 0 2s  Z���        �v  Z���v  h���0 0 3s  Z���        �v  Z���v  h���0 0 4s  Z���        �v  Z���v  h���0 0 5s  Z���        �v  Z���v  h���0 0 6s  Z���        �v  Z���v  h���0 0 7s  Z���        �v  Z���v  h���0 0 8s  Z���         �Y  ~���Y  o���X X             1     �b  ����b  }���0 0                  �o  ~���o  o���X X             4     �v  ����v  }���0 0                  �v  ����v  }���0 0                  �v  ����v  }���0 0                  �v  ����v  }���0 0                  ��  ~����  o���X X             4     ��  �����  }���0 0                  ��  �����  }���0 0                  ��  �����  }���0 0                  ��  �����  }���0 0                                	�+    ?   ����?   ����        6   �� 	 Cbusprobe(  ����E  ����  ����f  ����  	remainder     �7  ����7  ����Z Z 	remainder  ����         �^  ����^  ����0 0 0[  ����        �^  ����^  ����0 0 1[  ����        �^  ����^  ����0 0 2[  ����        �^  ����^  ����0 0 3[  ����                          H+       ����   �������{   n  ��  �����  �����  �����  ����  quotient     ��  �����  ����Z Z quotient�  ����         ��  �����  ����0 0 0�  ����        ��  �����  ����0 0 1�  ����        ��  �����  ����0 0 2�  ����        ��  �����  ����0 0 3�  ����                          H+       ����   ����         ��  CbusZ  ��  Csegment*  W���*  W����*  H���*  H����*  W���*  H���   5 �Z  �?  ����?  �����g  ����g  �����?  ����?  �����g  ����g  �����g  ����?  ���� +  L �Z  ��   %����   /�����   %����   %�����   /����   /��� _  u �Z  �  ����  ������   �����   �����  ����  ������   �����   ������   ����  ���� !  � �Z  ��   �����   ������   �����   ������   �����   ������   �����   ������   �����   ���� |  e �Z  ��   �����   ������   �����   ������   �����   ���� o  � �Z  ��   @����   @����R   B���R   $����R   $����   $�����   /����   $�����   /����   /�����   B���R   B�����   @����   B��� Y  � �Z  ��   @����   @�����   �����   ������   �����   ������   @����   ���� �  � �Z  �*  ����*  ������  ����*  �����*  ����*  ������  $����  ������   ����   �����   ����  �����  ����  $�����  $���o  $����o  J���o  $����o  J���o  J�����   ����   ��� � �   ��  Cnet0  �]  ����]  �����]  ����]  �����]  ����]  �����]  ����]  ���� A  � M�0  ��   �����   ������   �����   ������   �����   ������   �����   ���� �  � M�1  �2  X����   X�����   X����   X����2  ����2  �����2  ����2  X����2  ����2  �����2  ����  �����  ����  �����  ����  ���� X �  � �Z  �r  ����r  x����r  x���r  x����r  ����r  ���� C  � �Z  ��   �����   {�����   {����   {�����   �����   ���� �  � M�1  ��   &����   ?����H   &���H   &�����   ?����   ?�����   W����   ?�����   W����   W����H   &����   &���   � M�0  ��   r����   S����G   S���G   S�����   r����   r����G   S����   S���   � M�0  �G   ����G   ������   ����   ����G   ���G   ������   ���G   ���   � M�1  ��   �����   ������   �����   ������   �����   ������   �����   ����   � M�1  �G   ����G   �����a   ����a   �����a   ����G   �����a   ����a   ���� �  � M�0  �c  ���c  ����s  u���s  u����s  ���s  u����c  ���s  ���   � M�0  �a   ����a   �����a   ����a   �����a   ����H   �����H   ����H   ���� �    � M�0  �   }���   X����W   X���   X����W   X���W   X����   }���   }��� �  k �Z  ��  ~����  ~�����  �����  ������  �����  ������  �����  ~�����  �����  ����  �Z  �o  ~���o  ~����7  ����7  �����o  ����o  ~����7  ����o  �����7  ����7  ���� 	 �   testing               